
LIBRARY ieee  ; 
    USE ieee.NUMERIC_STD.all  ; 
    USE ieee.std_logic_1164.all  ; 
    use ieee.math_real.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity uart_comm_32_bit_tb is
  generic (runner_cfg : string);
end;

architecture vunit_simulation of uart_comm_32_bit_tb is

    --------------------------------------
    use work.uart_rx_pkg.all;
    use work.uart_tx_pkg.all;

    --------------------------------------
    package fpga_interconnect_pkg is new work.fpga_interconnect_generic_pkg 
        generic map(number_of_data_bits => 32,
                 number_of_address_bits => 16);

    --------------------------------------
    package uart_protocol_pkg is new work.serial_protocol_generic_pkg
    generic map(serial_rx_data_output_record => uart_rx_data_output_group
                ,serial_tx_data_input_record  => uart_tx_data_input_group
                ,serial_tx_data_output_record => uart_tx_data_output_group
                --------------------------------
                ,serial_rx_data_is_ready => uart_rx_data_is_ready
                --------------------------------
                ,get_serial_rx_data => get_uart_rx_data
                --------------------------------
                ,init_serial => init_uart
                --------------------------------
                ,transmit_8bit_data_package => transmit_8bit_data_package
                --------------------------------
                ,serial_tx_is_ready  => uart_tx_is_ready
                ,g_data_bit_width    => 32
                ,g_address_bit_width => 16
            );
    --------------------------------------

    use uart_protocol_pkg.all;
    use fpga_interconnect_pkg.all;

    package uart_protocol_test_pkg is new work.serial_protocol_generic_test_pkg
        generic map(uart_protocol_pkg);

    use uart_protocol_test_pkg.all;

    constant clock_period      : time    := 1 ns;
    constant simtime_in_clocks : integer := 15000;
    
    signal simulator_clock     : std_logic := '0';
    signal simulation_counter  : natural   := 0;
    -----------------------------------
    -- simulation specific signals ----

    signal uart_rx_data_in  : uart_rx_data_input_group := (number_of_clocks_per_bit => 24);
    signal uart_rx_data_out : uart_rx_data_output_group;

    signal uart_tx_data_in  : uart_tx_data_input_group   := init_uart_tx(24);
    signal uart_tx_data_out : uart_tx_data_output_group;
    signal uart_protocol    : serial_communcation_record := init_serial_communcation;

    signal number_of_registers_to_stream : integer range 0 to 2**23-1 := 0;
    signal stream_address : integer range 0 to 2**16-1 := 0;

    signal fpga_controlled_stream_requested : boolean := false;

    signal bus_to_communications   : fpga_interconnect_record := init_fpga_interconnect;
    signal bus_from_communications : fpga_interconnect_record := init_fpga_interconnect;

    constant g_clock_divider : integer := 24;

    signal uart_rx : std_logic := '1';
    signal uart_tx : std_logic;

    type std32_array is array (natural range <>) of std_logic_vector(31 downto 0);
    signal test_data : std32_array(1 to 5) := (others => (others => '1'));

    signal tuitui : std_logic_vector(31 downto 0) := (others => '0');

    signal transmit_counter : natural := 1;

    constant data_to_be_transmitted : std32_array :=(1 => x"acdcacdc", 2 => x"abcdabcd", 3=> x"12341234", 4=>  x"11111111", 5 => x"01010101");

begin

------------------------------------------------------------------------
    simtime : process
    begin
        test_runner_setup(runner, runner_cfg);
        wait for simtime_in_clocks*clock_period;
        check(data_to_be_transmitted = test_data, "words were not the same");
        test_runner_cleanup(runner); -- Simulation ends here
        wait;
    end process simtime;	

    simulator_clock <= not simulator_clock after clock_period/2.0;
------------------------------------------------------------------------

    test_uart : process(simulator_clock)
    begin
        if rising_edge(simulator_clock) then
            simulation_counter <= simulation_counter + 1;

            init_uart(uart_tx_data_in, g_clock_divider);
            set_number_of_clocks_per_bit(uart_rx_data_in, g_clock_divider);
            create_serial_protocol(uart_protocol, uart_rx_data_out, uart_tx_data_in, uart_tx_data_out);

            if transmit_is_ready(uart_protocol) or simulation_counter = 10 then
                transmit_counter <= transmit_counter + 1;
                if transmit_counter <= data_to_be_transmitted'high then
                    transmit_words_with_serial(uart_protocol, (0 => x"04", 1 => x"00", 2 => x"01", 3 => x"ac", 4 => x"dc", 5 => x"ab", 6 => x"ba"));
                elsif transmit_counter <= data_to_be_transmitted'high+1 then
                    transmit_words_with_serial(uart_protocol, read_frame(address => 1));
                end if;
            end if;

            if frame_has_been_received(uart_protocol) then
                if get_command(uart_protocol) = 2 then
                    transmit_words_with_serial(uart_protocol,write_frame(get_command_address(uart_protocol), test_data(3)));
                end if;
            end if;

            if simulation_counter = 8500 then
                    transmit_words_with_serial(uart_protocol,stream_frame(5));
            end if;


            init_bus(bus_to_communications);
            connect_data_to_address(bus_from_communications, bus_to_communications, 1, test_data(1));
            connect_data_to_address(bus_from_communications, bus_to_communications, 2, test_data(2));
            connect_data_to_address(bus_from_communications, bus_to_communications, 3, test_data(3));
            connect_data_to_address(bus_from_communications, bus_to_communications, 4, test_data(4));
            connect_data_to_address(bus_from_communications, bus_to_communications, 5, test_data(5));
            connect_data_to_address(bus_from_communications, bus_to_communications, 5, tuitui);

        end if; -- rising_edge
    end process test_uart;	
------------------------------------------------------------------------
    u_uart_rx : entity work.uart_rx
    port map(clock => simulator_clock   ,
          uart_rx_FPGA_in.uart_rx => uart_rx ,
    	  uart_rx_data_in  => uart_rx_data_in     ,
    	  uart_rx_data_out => uart_rx_data_out); 
------------------------------------------------------------------------
    u_uart_tx : entity work.uart_tx
        port map(clock => simulator_clock               ,
          uart_tx_fpga_out.uart_tx => uart_tx ,
    	  uart_tx_data_in => uart_tx_data_in  ,
    	  uart_tx_data_out => uart_tx_data_out);
------------------------------------------------------------------------
    communications_under_test : entity work.fpga_communications
    generic map(fpga_interconnect_pkg => fpga_interconnect_pkg
                -- , serial_protocol_pkg => work.uart_protocol_pkg)
               )
        port map(
            clock => simulator_clock                         ,
            uart_rx                 => uart_tx               ,
            uart_tx                 => uart_rx               ,
            bus_to_communications   => bus_to_communications ,
            bus_from_communications => bus_from_communications
        );
------------------------------------------------------------------------
end vunit_simulation;
